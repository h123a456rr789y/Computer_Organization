module Simple_Single_CPU( clk_i, rst_n );

//I/O port
input         clk_i;
input         rst_n;

//Internal Signles
wire	[31:0]instruction,regWriteData,readData1,readData2,Alu_result,Shifter_result,Alu_Shifter;
wire	RegWrite,AluSrc,Alu_overflow;
wire	[2:0]AluOp;
wire    [1:0] MemtoReg;
wire    [1:0] RegDst;
wire	[31:0]signExtend_tmp,zeroFilled_tmp;

wire    jump,Branch,BranchType,MemWrite,MemRead,Alu_zero;
wire    jr;
wire    [31:0]pc_now,pc_next,pc_end, pc_branch, pc_not_jump, pc_not_jumpReg;




assign jr = (instruction[31:26] == 6'b111111 && instruction[5:0] == 6'b001000) ? 1'b1 : 1'b0;


//modules
Program_Counter PC(
            .clk_i(clk_i),      
	    .rst_n(rst_n),     
	    .pc_in_i(pc_next) ,   
	    .pc_out_o(pc_now) 
	    );
	
Adder Adder1(					//PC+4
        .src1_i(pc_now),     
	.src2_i(32'd4),
	.sum_o(pc_end)    
	 );


Adder Adder_branch(  						//branch
		.src1_i(pc_end),
		.src2_i({signExtend_tmp[29:0], 2'b00}),
		.sum_o(pc_branch)
		);

Mux2to1 #(.size(32)) Mux_Jump(
        .data0_i(pc_not_jump),
        .data1_i({pc_end[31:28], instruction[25:0], 2'b00}),	//jump 
        .select_i(jump),
        .data_o(pc_not_jumpReg)
        );

Mux2to1 #(.size(32)) Mux_JumpReg(
        .data0_i(pc_not_jumpReg),
        .data1_i(readData1),
        .select_i(jr),
        .data_o(pc_next)
        );

Mux2to1 #(.size(32)) Mux_Branch(
        .data0_i(pc_end),
        .data1_i(pc_branch),
        .select_i(Branch & (Alu_zero ^ BranchType)),
        .data_o(pc_not_jump)
        );



	
Instr_Memory IM(
        .pc_addr_i(pc_now),  
	    .instr_o(instruction)    
	    );

wire [4:0]Reg_Write_addr;

Mux3to1 #(.size(5)) Mux_Reg_Write(
        .data0_i(instruction[20:16]),
        .data1_i(instruction[15:11]),
        .data2_i(5'b11111),
        .select_i(RegDst),
        .data_o(Reg_Write_addr)
        );	


Decoder Decoder(
        .instr_op_i(instruction[31:26]), 
        .RegWrite_o(RegWrite), 
        .ALUOp_o(AluOp),   
        .ALUSrc_o(AluSrc),   
        .RegDst_o(RegDst),
        .Branch_o(Branch),
        .BranchType_o(BranchType),
        .Jump_o(jump),
        .MemRead_o(MemRead),
        .MemWrite_o(MemWrite),
        .MemtoReg_o(MemtoReg)  
	);
		
Reg_File RF(
        .clk_i(clk_i),      
	.rst_n(rst_n) ,     
        .RSaddr_i(instruction[25:21]) ,  
        .RTaddr_i(instruction[20:16]) ,  
        .RDaddr_i(Reg_Write_addr) ,  
        .RDdata_i(regWriteData)  , 
        .RegWrite_i(RegWrite& ~jr),
        .RSdata_o(readData1) ,  
        .RTdata_o(readData2)   
        );


	


wire	[3:0]Alu_op;
wire	[1:0]FURslt;


Zero_Filled ZF(
        .data_i(instruction[15:0]),
        .data_o(zeroFilled_tmp)
        );

Sign_Extend SE(
        .data_i(instruction[15:0]),
        .data_o(signExtend_tmp)
        );

ALU_Ctrl AC(
        .funct_i(instruction[5:0]),   
        .ALUOp_i(AluOp),   
        .ALU_operation_o(Alu_op),
	.FURslt_o(FURslt)
        );



wire [31:0]Alu_input;	

		
ALU ALU(
	.aluSrc1(readData1),
	.aluSrc2(Alu_input),
	.ALU_operation_i(Alu_op),
	.result(Alu_result),
	.zero(Alu_zero),
	.overflow(Alu_overflow)
	    );

Mux2to1 #(.size(32)) Mux_ALU_Src(
        .data0_i(readData2),
        .data1_i(signExtend_tmp),
        .select_i(AluSrc),
        .data_o(Alu_input)
        );	

wire	[4:0]shift_tmp;
Mux2to1 #(.size(5)) Mux_Shift(
        .data0_i(instruction[10:6]),
        .data1_i(readData1),
        .select_i(Alu_op[1]),
        .data_o(shift_tmp)
        );

Mux3to1 #(.size(32)) Mux_FUR(
        .data0_i(Alu_result),
        .data1_i(Shifter_result),
        .data2_i(zeroFilled_tmp),
        .select_i(FURslt),
        .data_o(Alu_Shifter)
        ); 

Shifter shifter( 
		.result(Shifter_result), 
		.leftRight(Alu_op[0]),
		.shamt(shift_tmp),
		.sftSrc(Alu_input) 
		);

                     

wire [31:0] MemReadData;

Mux3to1 #(.size(32)) Mux_WB(
		.data0_i(Alu_Shifter),
		.data1_i(MemReadData),
		.data2_i(pc_end),
		.select_i(MemtoReg),
		.data_o(regWriteData)
		);		



Data_Memory DM(
                .clk_i(clk_i),
                .addr_i(Alu_result),
                .data_i(readData2),
                .MemRead_i(MemRead),
                .MemWrite_i(MemWrite),
                .data_o(MemReadData)
                );
              


endmodule




